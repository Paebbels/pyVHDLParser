use lib0.pkg0.all;

use lib1.pkg1.all ;

use lib2.pkg2.all; -- comment

use		lib3.pkg3.all		;

use lib4.pkg4.const4;
