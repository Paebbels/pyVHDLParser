entity/* comment0 */myEntity1/* comment1 */is/* comment2 */end/* comment3 */;/* comment4 */
entity /* comment0 */ myEntity1 /* comment1 */ is /* comment2 */ end /* comment3 */ ; /* comment4 */
