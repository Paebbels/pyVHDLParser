architecture rtl of myEntity is
begin
	process(all)
	begin
	end process;

	process(Clock)
	begin
	end process;

	process(Clock) begin
	end process;

	process(Clock)begin
	end process;
	
	process (Clock, Reset)
	begin
	end process;

	process(Clock) is
	begin
	end process;

	process(Clock) is begin
	end process;

	-- proc:process(Clock)
	-- begin
	-- end process;

	-- proc: process(Clock)
	-- begin
	-- end process;

	-- proc : process(Clock)
	-- begin
	-- end process;
end architecture;
