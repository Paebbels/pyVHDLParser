package
body
myPackage0
is
end
;

package    -- comment0
body       -- comment1
myPackage1 -- comment2
is         -- comment3
end        -- comment4
;          -- comment5

package-- comment0
body-- comment1
myPackage2-- comment2
is-- comment3
end-- comment4
;-- comment5

package    /* comment0 */
body       /* comment1 */
myPackage1 /* comment2 */
is         /* comment3 */
end        /* comment4 */
;          /* comment5 */

package/* comment0 */
body/* comment1 */
myPackage4/* comment2 */
is/* comment3 */
end/* comment4 */
;/* comment5 */

package body myPackage5 is end;
package body myPackage6 is end package body;
package body myPackage7 is end myPackage7;
package body myPackage8 is end package body myPackage8;
package body myPackage9 is end package body myPackage9 ;

package body	myPackage10	is	end;
package body	myPackage11	is	end	package body;
package body	myPackage12	is	end	myPackage12;
package body	myPackage13	is	end	package body	myPackage13;
package body	myPackage14	is	end	package body	myPackage14 ;

package body myPackage15 is 
end;

package body myPackage16 is
end ;

package body myPackage17 is
end package body;

package body myPackage18 is
end package body ;

package body myPackage19 is
end myPackage19;

package body myPackage20 is
end myPackage20 ;

package body myPackage21 is
end package body myPackage22;

package body myPackage23 is
end package body myPackage23 ;

package body/* comment0 */myPackage24/* comment1 */is/* comment2 */end/* comment3 */;/* comment4 */

package body /* comment0 */ myPackage25 /* comment1 */ is /* comment2 */ end /* comment3 */ ; /* comment4 */
