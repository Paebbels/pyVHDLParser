package
myPackage0
is
end
;

package    -- comment0
myPackage1 -- comment1
is         -- comment2
end        -- comment3
;          -- comment4

package-- comment0
myPackage2-- comment1
is-- comment2
end-- comment3
;-- comment4

package    /* comment0 */
myPackage1 /* comment1 */
is         /* comment2 */
end        /* comment3 */
;          /* comment4 */

package/* comment0 */
myPackage4/* comment1 */
is/* comment2 */
end/* comment3 */
;/* comment4 */

package myPackage5 is end;
package myPackage6 is end package;
package myPackage7 is end myPackage7;
package myPackage8 is end package myPackage8;
package myPackage9 is end package myPackage9 ;

package	myPackage10	is	end;
package	myPackage11	is	end	package;
package	myPackage12	is	end	myPackage12;
package	myPackage13	is	end	package	myPackage13;
package	myPackage14	is	end	package	myPackage14 ;

package myPackage15 is 
end;

package myPackage16 is
end ;

package myPackage17 is
end package;

package myPackage18 is
end package ;

package myPackage19 is
end myPackage19;

package myPackage20 is
end myPackage20 ;

package myPackage21 is
end package myPackage22;

package myPackage23 is
end package myPackage23 ;

package/* comment0 */myPackage24/* comment1 */is/* comment2 */end/* comment3 */;/* comment4 */

package /* comment0 */ myPackage25 /* comment1 */ is /* comment2 */ end /* comment3 */ ; /* comment4 */
