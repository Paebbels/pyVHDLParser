context OSVVM is
	use OSVVM.Scoreboard.all;
end context;

context
	OSVVM
		is
			use OSVVM.Scoreboard.all;
				end
					context
						;

context OSVVM is use OSVVM.Scoreboard.all; end context;
