use lib0.pkg0.all;

use lib1.pkg1.all ;

use lib2.pkg2.all; -- comment

use		lib3.pkg3.all		;

use lib4.pkg4.const4;

use lib5 . pkg5 . const5;

use
lib61
.
pkg61
.
const61
;

use
	lib62
		.
			pkg62
				.
					const62
						;

use lib7.pkg7.const71,lib7.pkg7.const72;

use lib8.pkg8.const81, lib8.pkg8.const82;

use lib9.pkg9.const91 , lib9.pkg9.const92;
