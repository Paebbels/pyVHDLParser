package pkg0 is
	function func0 return integer;
end package;

package body pkg0 is
	function func0 return integer is
	begin
	end function;
end package body;
