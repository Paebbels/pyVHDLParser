architecture rtl of myEntity is
begin
	process(Clock) is
	begin
	end process;

	process(Clock) is begin
	end process;
end architecture;
