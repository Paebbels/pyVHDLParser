package pkg0 is
	function func0(a : integer) return integer;
end package;

package body pkg0 is
	function func0(a : integer; b : integer) return integer is
	begin
	end function func0;
end package body;
