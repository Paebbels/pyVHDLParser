library library0;

library library1 ;

library
	library2
		;

library 
	library3 
		; 

library library4;  -- comment

library -- comment1
	library5  -- comment2
; -- comment3

library-- comment
	library6--
	;-- 

library
library7
;

library library81, library82;

library library91, library92;

library
	library101,
	library102;
