entity
myEntity0
is
end
;

entity    -- comment0
myEntity1 -- comment1
is        -- comment2
end       -- comment3
;         -- comment4

entity-- comment0
myEntity2-- comment1
is-- comment2
end-- comment3
;-- comment4

entity    /* comment0 */
myEntity1 /* comment1 */
is        /* comment2 */
end       /* comment3 */
;         /* comment4 */

entity/* comment0 */
myEntity4/* comment1 */
is/* comment2 */
end/* comment3 */
;/* comment4 */

entity myEntity5 is end;
entity myEntity6 is end entity;
entity myEntity7 is end myEntity7;
entity myEntity8 is end entity myEntity8;
entity myEntity9 is end entity myEntity9 ;

entity	myEntity10	is	end;
entity	myEntity11	is	end	entity;
entity	myEntity12	is	end	myEntity12;
entity	myEntity13	is	end	entity	myEntity13;
entity	myEntity14	is	end	entity	myEntity14 ;

entity myEntity15 is 
end;

entity myEntity16 is
end ;

entity myEntity17 is
end entity;

entity myEntity18 is
end entity ;

entity myEntity19 is
end myEntity19;

entity myEntity20 is
end myEntity20 ;

entity myEntity21 is
end entity myEntity22;

entity myEntity23 is
end entity myEntity23 ;

entity/* comment0 */myEntity24/* comment1 */is/* comment2 */end/* comment3 */;/* comment4 */

entity /* comment0 */ myEntity25 /* comment1 */ is /* comment2 */ end /* comment3 */ ; /* comment4 */
