
entity    /* comment0 */
myEntity1 /* comment1 */
is        /* comment2 */
end       /* comment3 */
;         /* comment4 */

entity/* comment0 */
myEntity4/* comment1 */
is/* comment2 */
end/* comment3 */
;/* comment4 */

architecture    /* comment0 */
rtl3            /* comment1 */
of              /* comment2 */
myEntity3       /* comment3 */
is              /* comment4 */
begin           /* comment5 */
end             /* comment6 */
;               /* comment7 */

architecture/* comment0 */
rtl4/* comment1 */
of/* comment2 */
myEntity4/* comment3 */
is/* comment4 */
begin/* comment5 */
end/* comment6 */
;/* comment7 */
