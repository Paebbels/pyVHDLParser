architecture
rtl0
of
myEntity0
is
begin
end
;

architecture 
rtl00 
of 
myEntity00 
is 
begin 
end 
; 

 architecture
 rtl000
 of
 myEntity000
 is
 begin
 end
 ;
