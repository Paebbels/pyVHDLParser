architecture
rtl0
of
myEntity0
is
begin
end
;

architecture 
rtl00 
of 
myEntity00 
is 
begin 
end 
; 

 architecture
 rtl000
 of
 myEntity000
 is
 begin
 end
 ;

architecture    -- comment0
rtl1            -- comment1
of              -- comment2
myEntity1       -- comment3
is              -- comment4
begin           -- comment5
end             -- comment6
;               -- comment7

architecture-- comment0
rtl2-- comment1
of-- comment2
myEntity2-- comment3
is-- comment4
begin-- comment5
end-- comment6
;-- comment7

architecture    /* comment0 */
rtl3            /* comment1 */
of              /* comment2 */
myEntity3       /* comment3 */
is              /* comment4 */
begin           /* comment5 */
end             /* comment6 */
;               /* comment7 */

architecture/* comment0 */
rtl4/* comment1 */
of/* comment2 */
myEntity4/* comment3 */
is/* comment4 */
begin/* comment5 */
end/* comment6 */
;/* comment7 */

architecture rtl5 of myEntity5 is begin end;
architecture rtl6 of myEntity6 is begin end architecture;
architecture rtl7 of myEntity7 is begin end rtl7;
architecture rtl8 of myEntity8 is begin end architecture rtl8;
architecture rtl9 of myEntity9 is begin end architecture rtl9 ;

architecture	rtl10	of	myEntity10	is	begin	end;
architecture	rtl11	of	myEntity11	is	begin	end	architecture;
architecture	rtl12	of	myEntity12	is	begin	end	rtl12;
architecture	rtl13	of	myEntity13	is	begin	end	architecture	rtl13;
architecture	rtl14	of	myEntity14	is	begin	end	architecture	rtl14 ;

architecture rtl15 of myEntity15 is 
begin
end;

architecture rtl16 of myEntity16 is
begin
end ;

architecture rtl17 of myEntity17 is
begin
end architecture;

architecture rtl18 of myEntity18 is
begin
end architecture ;

architecture rtl19 of myEntity19 is
begin
end rtl19;

architecture rtl20 of myEntity20 is
begin
end rtl20 ;

architecture rtl21 of myEntity21 is
begin
end architecture rtl21;

architecture rtl23 of myEntity23 is
begin
end architecture rtl23 ;

architecture/* comment0 */rtl24/* comment1 */of/* comment2 */myEntity24/* comment3 */is/* comment4 */begin/* comment5 */end/* comment6 */;/* comment7 */
architecture /* comment0 */ rtl25 /* comment1 */ of /* comment2 */ myEntity25 /* comment3 */ is /* comment4 */ begin /* comment5 */ end /* comment6 */ ; /* comment7 */
