package body pkg0 is
	function func0 return integer is
		constant const3 : integer := 15;

		/*function func1 return integer is
			constant const4 : integer := 20;
		begin
		end function func0;*/
	begin
	end function func0;
end package body;