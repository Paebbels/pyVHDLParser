architecture
rtl0
of
myEntity0
is
end
;

architecture 
rtl00 
of 
myEntity00 
is 
end 
; 

 architecture
 rtl000
 of
 myEntity000
 is
 end
 ;

architecture    -- comment0
rtl1            -- comment1
of              -- comment2
myEntity1       -- comment3
is              -- comment4
end             -- comment5
;               -- comment6

architecture-- comment0
rtl2-- comment1
of-- comment2
myEntity2-- comment3
is-- comment4
end-- comment5
;-- comment6

architecture    /* comment0 */
rtl3            /* comment1 */
of              /* comment2 */
myEntity3       /* comment3 */
is              /* comment4 */
end             /* comment5 */
;               /* comment6 */

architecture/* comment0 */
rtl4/* comment1 */
of/* comment2 */
myEntity4/* comment3 */
is/* comment4 */
end/* comment5 */
;/* comment6 */

architecture rtl5 of myEntity5 is end;
architecture rtl6 of myEntity6 is end architecture;
architecture rtl7 of myEntity7 is end rtl7;
architecture rtl8 of myEntity8 is end architecture rtl8;
architecture rtl9 of myEntity9 is end architecture rtl9 ;

architecture	rtl10	of	myEntity10	is	end;
architecture	rtl11	of	myEntity11	is	end	architecture;
architecture	rtl12	of	myEntity12	is	end	rtl12;
architecture	rtl13	of	myEntity13	is	end	architecture	rtl13;
architecture	rtl14	of	myEntity14	is	end	architecture	rtl14 ;

architecture rtl15 of myEntity15 is 
end;

architecture rtl16 of myEntity16 is
end ;

architecture rtl17 of myEntity17 is
end architecture;

architecture rtl18 of myEntity18 is
end architecture ;

architecture rtl19 of myEntity19 is
end rtl19;

architecture rtl20 of myEntity20 is
end rtl20 ;

architecture rtl21 of myEntity21 is
end architecture rtl21;

architecture rtl23 of myEntity23 is
end architecture rtl23 ;
