architecture arch of ent is
begin
	assert False report sdfjcsdfcsdj;
	assert False report sdfjcsdfcsdj severity note;
end architecture;
