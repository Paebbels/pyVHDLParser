package pkg0 is
end package;

package body pkg0 is
end package body;
